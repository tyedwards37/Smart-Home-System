PK   0!�S��!01  ��    cirkitFile.json�}ێ�ȑ�����߽��V��I,�����P)�6+K�AC�?�ߴtFFUF8��,;6j���]���C���_��y��<��q���������[2�7���^�����pw�{z���������?�?����0��q�����f����;(C�W.�A%���gsH:��N������z�������Q=vw��><����cj������O����]t�Cg�U�wF9���ՠ����>���A��Rp�ΰ9��ױQB�a���+����"�csp�/�~�=��ϖ���w�́��w�́��w��!1�2��%�q�ڧ�|�T�9)��IeGN��c���wޱ�N�ݙ�����+ x2L���}�;=6�Ă���!ty�l�kV�@��o�gE�<�d>�bCL,��bb�����#�R����V�c��e�T�6*=dM�$c�l��,E�����R������߭�_��]ڛ�k��H"ײȶ�7���5�ߑ�_���y|�}|~a��5�������������3�W?@�> ?J�!��"���I�`��Ȱb#�� ��g���e�B�P�jddh���e�B�P������e�B�7��O��b!�`�y��F�i����B���͂?�b�1bb�<�~�����e�i8.�Ă�{�!&�^�1���%l��`z�1���N��v�n���n-�l��������Z������;��w�I^��u�����i��1����K�~_�X��6�.��,�}����������gCL,�~�1�`-�q�a\:ޞ�t��wwui0��,������&o�|��ᬶ'�M���/!��yk]΃N�RM�"C�20���"�{3�G�G���*m`p�7g���V��}mf��m�g"�;�T��!ޙE�;��#,;²��V�v��a�MQ+V;��ʎ����]�jeGXvz��E�vPv�ew���]B�V��KC���g�I���g��B��]ف�������_����u����mK`�� ���_�p���`��_�*���`��_�C�9�R�T�~<D~p�C�tˏ���f@�~��ˏ���6F�~�Ԁ��̯l��N^��̯l���g������M�`�������]�`�������m�`�������}�`���������`�������}�`�������m�`�������]�`�������M�`�������o3���.����B~<Zx<�\��ł�,?�+;�����,?�wV3?W����f�f��ǂ��˭����]��}<Zx<�\��ɂ�',?�+������',?�+�����',?�+�����',?�+5����',?�+�)��9�������`�������� `�������Z&`�������*,`��{dЛd���e��Q��3N_����A��/��`��_)����`���y��~�-7����x��xL��ُg?X~�W�)a����ˏ��J%(�~��ˏ��J+�~��ˏ��J�-�~��ˏ��J�0�~��ˏ��J�3�~�*�2��Ń�N_��̯T��N_��̯����}��#0�R��8���#0�RW�_ �X~�W����X~�w^S��+U;�d&S.p�R?�K��e�.K�nl~Y@sc���[k��_��Za��������ey76������e1ۭf�5;��U�omϴ��X�홶W���=���k��g�_u����\�Ǵ��Lέ��W�
��=���3��g�_u"�֎�iG�m�^�⽕
������>�twcX����[�����u�Ƚ}fݞ��c��Wo�}ŗ'm���Ъ󰶶����:�j{!�%��pn����8�O��{�w�2Ӎ\$���-����ļ�e�������_��u�z�2�ꤠ�홁pu:����.�:�f� 3�Np�ڞi��i���o� ��������"��"��"��"��"��"��"w�i�i�i�i�i�i�i�i�i�i�;ϴ�Ĵ�̴�̴�̴�̴�̴��n���ʑ�q��N�{�h��$����`�+�oM���}6vԽ�v����u�vP>Y�6i����75_�;�G�
�#��*��SC6���{��M������qԪ��+�QV���<`�p�)MO���gSs���;����bo��Q����j^������v��l��{�ٛ��?{S��goj���f��A���q��c>(o��ޘnԯ<{S�W�{���T[��yzqY;�m�~��)�dl�w�����6ݝ=R�6��twý��Y�ݹ���$Mw��2\���xw�$��I���s�sw����`��y���$���qQ�Yކ��V'��n��v�Skm�纻ՉŶۋM��ݞ=��rx��x�����tS�B�r���1�AO����χ��˯={���fϹ9��׾��߇~�)�rc0�sdUߏ�9"3�)��vM��C��毄�}OS���ޥ���Ѩdz��}��{k\�_ˆ�����:��==솇��7o�L�L�n����������h�1�@@��t�#�{��#�b�%��0z���ȣ��t��1�@@���F  ]bi����<;�R�2�(�洏H�~�]x���	�a~�`�����	�	漏H{���#$2�9p���8�|8��8
Iϛ	@�2�g10?n`ѷ���y瘜p����{�ݷLN0?~B��뙜`~���I&|����'�o~��������;���������	)���w��G$��������i�&���a~����[,̏�޽������7��J��>�������X�G!�yc�,�0?�B��('X<na~���Z�AL���l�8��U̏������	7&�!�y�l\����i

�6LN0?~B��&O����6:�`~���z����0?�B��>'��0?�B���C'����MX<�a~��罓 N�x���8
iޜ]�~p�}CLN0?`~<��U��}�u��`~<<��h"�ӊ�^�Ⲛ�R��B���-����j�|h�+_��*�]/k=bt��"t]��W�|#F��"�]k�]�����JG�q%�$�uʻDt��Y�Q@�+�p�� ]/k�c��J"\�ED���$��W���zG�*��D���e5|8*0��J�\�
\Vɇ��U�+�p-k�E�%�,�dؒ۲�YF[�L�dؒ۲F[F[�l�dؒ۲�\F[��K�-ɰ-k�e����Dؒ۲�_f�K&[`��Ej+���L&&dؖ�2��dc"lI�m�S"��D�C2lI�m�#��LV&dؖ=>"���L�-ɰ-{�d����Dؒ۲�JF[��L�-ɰ-{�d����Dؒ۲NF[��L�-ɰ-{�d����Dؒ۲'QF[��L�-ɰ-{+e����Dؒ۲GTF[��L�-ɰ-{]e����Dؒ۲gWfa��
E��� �L^fe�2�$ö졖�V&/aK2l�^p�y+�ZQh��L^fe�2��� ��L^�� �L^fe�2�$ö���V&/aK2lK�me�2�$ö�|��V&/aK2lK�
me�2�$ö�����̗��%������2y�[�a[j��h+����%������2y�[�a[j��h+��Lh+�L^�d�1:��l�-��L^�d�2�$ö�>��V&/aK2lK'mev����e� d�2'����%������^&/aK2lKm0me�2�$ö�8��V&/aK2lK�6me�2�$öԜ��V&/aK2lK�<m��|����˼L^�e�2�$ö�2��V&/aK2lKMFme��Dؒ�R[RF[��L�-ɰ-52E�2y�[�a[j}�h+����%��f���2E��2�K�/gD�S��O*朔�뤲#�|Ї1��R�k:oDY�M�e���F��:�QV*ooDY���e���F��z�QV*HoDY�����@Ƌ�޵C_��`�w�֭0^;�t+Ɔ׎	�
���c=�|0Ɗ�λ�
���S%��`�x��ƭ0+^;!qk�����9��1�VP(�lŗg�n����>Fv+̳_���f����֭0�y���y�[a0V�v��֨o�`�0_�v��VPD���k'�m�9�����0���sl�9Zqu�V�g+�<�kk��lŗǚm�Y9�u+Ɗ��g�
3[�R��`�x�ࢭ0��b�x��0_�v��V�/^;�f+Ɗ���ƊƊƊƊ#Ɗ#Ɗ#Ɗ#Ɗ#Ɗ#Ɗ#h�c�c�c�	c�	c�	c�	c�	c�	c�	c�	4Z��ℱ⌱⌱⌱⌱⌱�|Պs7��٨t:��U��+�l>ꆃ5�g��P����gcG�+m�^��u�vP>Y�6i��:�&��\HG=j�TH)�V�����|<�x�u.M(W��C0}��b��u�U��2#�CLiz����&���R��/�{}�*�^O����~�^�8��Ҙ��w�uiB��K�U]�P��b�0���]�:7�<��&�����F}]�&���ҧ�h��1Oo:k��-�bȚ�I�Fڭ����6�<����ݻ(��XM���⯍7�́�������s�����&�9��Τ��;�s����D�Y�����`N3-��	m0���F�ՙ�6�$O����A�\e7*��(���z��6Y[��C��:�ЄB��C���Di��>S0�G��`T�Ȫ��sDf�n���&��>�	�z���4�aZ�]:LqY4*�ިa����冈�	���u��==�>>uO��۟��n?���?==v�_��~V7��C���l	F  =��F  =��F  =G	F  =GF  =G/F  =GBF  =GUF  }��0.�qn�	�QH��b8�|7��7
ICd'��&�G!��U'�'�G!��bZ'�70?�B��e�N��������q�>�f�p��q��($}\g������QH���	��̏���qm:&��q��($}\5��I�������q�>n�p��q��($}ܶ������QH����	��̏���q��̏;�G!��&'ܘ8nP��̏���q��̏;�G!��. '�w0?�B���I����0?�B�ǝSN0?�a~���{�0�p����M��0?�B�ǭkN0?�a~�����0�`~<��8
I��a8��x���5�핯��jh�c�* *�p%�zWUUC�u��J"\�����F�*��D��]U��
�U�+�p��.]��$���)ѵ*nQ@�+�p�b]���$��W���Z�Q��Jp%�zWU�F�u��J"\���f�F�*��D��5�2��L�%dؖ��2�
e]Bi�L�E2��d^"lI�mYk.��L�%dؖ5�2��d`"lI�mY�/��L&dؖ=2��db"lI�mً!��L6&dؖ=%2��dd"lI�m�#��LV&dؖ=>22y�[�a[�*�h+����%�eϕ��B3bBSb2y���ˌL^&dؖ=p2���e"lI�m��'��L^&dؖ=�2���e"lI�m�[)��L^&dؖ=�2���e"lI�m��*��L^&dؖ=�2�d�2�$ö�=��V&/aK2l�jme�2�$ö���Vh���rE�����eV&/aK2l��|me�2�$ö���V&/aK2lK�me�2�$ö�|��V&/aK2lK�
me�2�$ö������e"lI�m�%"��L^&dؖ�(2���e"lI�m��"��L^&dؖ52�
�$�J&��9�����e"lI�m�$��L^&dؖ�G2���e"lI�m��$��L^&dؖZT2���e"lI�m��%�����Dؒ�RLF[��L�-ɰ-5�d����Dؒ�R�MF[��L�-ɰ-5�d����Dؒ�R;OF[�*Be>d�2/��y��L�-ɰ-�e����Dؒ�R�QF[��L�-ɰ-�%e����Dؒ�R#SD� ����%��֧��2y�[�a[j��h+�����6�_��ާ�|�T�9)��IeGN��c�����aވ�R�v#�J5ٍ(+u�7��T�ވ�R+{#�Ju�(+��7��T�ވ�R�y�Ձ�c�k��n�����Ѫ[a0�v��V���c�k�qn��`���R�c�kgAn��X�ډ�[a0V�v���^c�k�n��+^;Vo+Ɗ���
���#��`�x� ��0+^;�l+("�X��9`[a0V�v��V���i�5��X���Q[a0V�v>�VPb��ⵃ���`�x�x��0+^;�g+Ɗ׎��
��‱� ��Xq�Xq�Xq�Xq�Xq�Xq�Xq�Xq�Xq�Xq�a�8b�8b�8a�8a�8a�8a�8a�8a�8a�8�F�1V�0V�1V�1V�1V�1V�1V��Zq�;:��C���J4xe��C�p����T����l�{���+�Nu��'kB�&>_�҄r��G�
�#��*��SC6����Υ	�*w���V]^����tPf�p�)M��0s؄��r�SjB��%bo��Q����8xՏ���Y����.M(WuiB��K�U]��!t�2�+V���|P�d��1ݨ��҄r�^�4�m�>��Mg�T��QYS2��H�ۂ��r�v[P���&���@��>�	�j ӄr5�iB��4�\�bڬd��>�������m0W-8N����zg��~P��Yz���>��^�	��{jB����~�}�`��ʍ��ΑU}?���\�&��OԄr�o�{��0��.��,�Lo԰�~o��rCDՄ���z;��?톇������߼5���/w���݇��0�ww������x�����t����a�yןn��P�X5����#�5�̅.��8�K�Pf�D���8;^��=�&�N��MFroO�IL��}�M~2maB`���q.Ϥs��K'�悹���m��i�4[9��慣�ۯ��֠�{��ؚpooy	�����qo��gwf��4��ܻ�8�Ɯ�{�ĸ;3(%�Yc/̻[��c�;��wlwg9���,�۱��qvl_�bt��,��5:��X�:��j{�Kи�0SB���k�W��q�ЫuŹP�պR](�j]�u��s�}�W����3Z`��o͂;�x��b��E���3�n�C7zǱL�v��x����9tuy:�O?�f.�?=�y�����,Ə�_���O�͏���C����/O#.#�T�b����/'F����˚O�L+aXpg� ,ؓLk���)|��
=�aŝ�°�N�������߿�< �{:Â;+�a��İ��bXp�
1,�3�̉C	��!�sC�9�!��TĐ`�-bH0�1$�3��	ǿI��|Ѽ�JLL̛�����"S4^l����g4E���M�x�y~S��9��l�h�<���_7�)A �@E#���_��x�2�˝g��2L�b��ge'Z7�Ow���O��x������vO�Ow���?s^u�!���콽�����I���-�L���|g;)�'ņ��Nr&W[�����t&)6��7�3Y�!��1�ɂ���L����T�3�c�+E ?L�#>����\1|1Cpy �/0��m. <c\�� ������< n� ~����G,py�q��bS�b�LZ _<c\�b�Q�x��V'3N6 O=c\�
LZ �mj�M�I�M����1.h��=}<�K+�a(��5 �n�mf�k ^�,�L/o^��^�0��xy[{y������hb8�����-�������� /����3j�< ��q>�>������-�S�1��\3C��� �~8���c��QC\��g��3C;��f�O�������:��uu�L�������f�L}��1��)�
�{�/�c��yW\ _������'nqy |�G��b[p�|}<4���z�{�c��e.��N��;[p�aa3���f��t��U� h�!�h��ɿ������e[�f�R�j�Lu�uu��V�^W���V��Vt��+��T�\�]�b`��3խ�2յP~gx ~�G`~S�ρ���#0�)�����a���p��`����O�"X��ˏ���V�C�K�wǆ���t���|��3��ˏ���*U���M͐�˒Z��ؔ��	Ͱ,Fk��	͐��Rf����̐��2l���̐���o�/���c$E'-`�e�;�,�y�!����hѹ�!��}h�	��a�#������a���Р�0CB3,�O���0CB3,[e���0CB3,�z���0CB3,�����0CB3,;����0CB3,ۻ���0CB3,{����0CB3,����0CB3,�����0CB3</m�Y.re�a��!4aZ �U ��Xt�fHh�e�'ZCt�fHh�uE��w���1������b.띾���+@'55a��Ƣ�0CB3,�����0CB3,����0CB3,�����0CB3,����0CB3,���:���!��Bh�Y�!��"
h�Y�!��h�i�!���h�Z�Z�y��y��W���c$E�-`��h�,�i�!��
'h�i�!������ʞ���&L��
����b�	Ͱ��k��Y�!��>h�Y�!���Ch�Y�!���Ih�Y�!���Oh�Y�!���Uh�������i�G�-����a)������a)s��=�fHh��DZCt�fHh���XÀ�S�	Ͱ�Ck��S�	ͰT�Ckx���cB��g�OU��Dnl__�ؾ�����df��B��Si����W�T7��*�nl_�*�j?l�Z`}|�V �և�m�Za}�V ��Ǿm�Zb}:�V �/�Zb}6�V �%��}m�Zb}��V �%��Rm�Ӹ��pN�yAԭx�^�V�Ώ܊�pR���-18x�\D�¡n��ǵ��4��q�Bmq���:���� �P��|�cc��f�9��©*��Y-������������r���v��V<���{lX8|.s�&_���oԇPl������� \�[���k���|{$�k��k��k��k��k��k��k��k��k��k��=(ŵ�ȵ�ȵ�ĵ�ĵ�ĵ�ĵ�ĵ�ĵ�ĵ���Zb�Zb�Zb�Zb�Zb�Zb�Zb~�s7��٨t:��U��+�l>ꆃ5�͓4���>;�^i;�ʅ�S]���ɚ��I�ϯݿ��+�'��}R!u���Z%�wjȦ��`�ap�ݿ��+�w�`�8j�����(��@eF
����0��S5�����O���+_�!�&�U�����U?N/qlgi���מ���+������oj���!C�ezW��*����ɾ?xc�Q���M�_{�}�>Zm�>���e�T��s��d���vufoVF������&���:�2n�W�֮;4�-��+C}Mp�X��Xh\=�eVƀ��FjW�����/Z/i�[�J3^�b}�w�6߆Wk�mx��mx��O��1V��89�n
QT�QN�A�:f5�ɗk��|���^�6������h�[8�s�a�~�}�謏ʍ��ΑU}?��:���4���ij�Z��4u�Z�]:L!^4*�ިa�����WC���G������n�{z�M�o��|�i߼����b&�ek._Hy��K.ޡx�����y�}6�����i�F��&������Jg�<������َ�.t����e[Z�G=ؙNiaK[Z�������+-\i�J7?Ai�JWZ�����/-|i�K??ti�K_Z�����E(-BiJ�0�TZ��"�����E,-biK�XZ��"�Җ����E*-Ri�J�TZ��"���H��(-Ri�K�\Z��"��������7�9_^�Ԡ%19kВI�5h	�k���Ĭ�[��s�~���Tl��<��Ԩ�=U�Z|�%&����N�ǧ�Mvӏ̅������/�X�ZCQ��3v��f�J[�����g3�gc�����D��Y�U�
ߺ�f���Y]�(�z��|u֪��Q�2���O��(2y�<��Ԍ��fU0�+$�3��g2�؇X1$�e�Y���q� �\1S3���b� ]�Q�̧c��W�k���{Xcekc�kJ���uT�X�㰖d�����r���p�H���E��V8��Z���e��/9bnwʚ�X�@��dͱ,i��y�h��n߹�z�q&��E,���+-��dv��GD�O��+-���t�~a,ð�ʗ��BNO˙�X҂��ZV?˴[{%�3�n�r�]����Q��q{af�{-�5�NY�X���J���s��h���Zn��N/G��W?����{����2l�/��y{����W��/~�矨��<�d���O���=�����O��)<����O��)=�����O���NjP-}��փNzP-��Z:)B�$t��jM�	բ�I�U��*T�B'Y��Ŝt1�.椋�u1���Ŝt1�.椋�u1']L��9�bj]�IS�bN��Zs��Ժؓ.��Şt��g����w/�����a����SqM�x�;����qgޜ�)�õߏ����3��ى��{*ӌ?��?>��Ow�<�����?ŝMB||z��/�"�ݟʟ˯�7��*���b�&�t7ѽ������/��M�7o�����������>������8��Ow�������{�O���C7<}z_#��L���� L&*��{�{�t�Q�C1N���O��6���/��I�B��'��q�B7z���z�s�"�����{G�<pw���m��7��<<�M��;���a����qx?>��ɛ7�6���������_�s���������4��Cf�ϟߞ~pk-�J:�<�{�k[p^z��w痛~0gO������}q�	���ܺ!�7/u��Z.]��./�^��U_,`���X��2��jM�.S���6f
G�.�N�w� k�Er�Ew~�
\u�2Z:o��
\}�2�����e���v���.]����
Z���B�?G˶��ڲ��/oz��T4+?�xy�������&��@-bX�K�k7�tՂ�Z��vrKW�.r��������ڵ︖h-����mRaft�G���]��eX�M�/��L���j0��l�̷1[��m̖.��R���j���l�
,Q���j0��l�̵1[���m̖.��b���j���l�
,��[�e���j0:�eZ[���~��=F��5_�3��rY��偳=��.^Uc�!ŉ�|UX�Z�jk2��l<ED+XWM1�y�>�����9�?͉��~��i��o���cNDo����/���?�s�����S�?'�/.��Z�y��9����"�,9�e9���������KG��x�Ι� ��ޏ��|&�����a��/��?�l�CI?�]ߘ����?�g��������G�Oe`!'�2�_�S?>��_�����|���/X��t�S�t���ە���M�M�O�;ih�˜;�!z��nJ�����W#كsqH��.s�5�9������T���/��dK,7��/:���;�`?�Ӗ&����r��y�
[d5�5��m���"��t%�U���gw!�������3u�.�7ƥl�)��C��7��i���<�(t�w ��-����׊&}~	#���=��ݧ{�кI����9���N�e������Pg;������U��N&v1�Ύ�xi3M۴F�� ���_��6b��l�;=��e���ҳ���y����a�9�r��1��_�n1�������o��^OQ�� +�������c�7D��٬�d�ּ�N�t�s/-q0�}�Ք���V�'R��Nn����Us<M��,qvI/Ɇe{sɴ]�W-���_�lq[�h	^�}wx�t�����*mƏs���T�1�Z_,0�d�)��b�{�7�f��<�,��I�������`���TF�c,fz��}M��ɥ���mf�}�wa2e�LO���"ݒ�:Ѳ8�>�|��l�{P��J*Ȩ�}���]�$#��D[6_Z�s�yn;e2�v�(�S&/Gvr|����2����\\��9��>��֠Lc�P�t���w/�޿��yĮ���S���C:^t��ӸՅ�]���:�]w1�3��.f\U��sQ�r����oN�x��Ϻ-���p[�v!��E#�f��4��M���S�k��Ôx�7*�N�q�d헦ݴi��)���[=��L��}��j?�/�����8R�^\'�*��������-��{؏'_9��{ɒjx��i|}r����G���笃C��4��LY��rɪ���:�)T3C��\���AS��o��=>U���cS�Ő���돿~���E�c��o2Ts��s�\���d�:D�XMS�����#�[w19���/�ֻ�4?���PK   0!�S��!01  ��            ��    cirkitFile.jsonPK      =   ]1    